// config.sv: Basic configuration file

// Define address width and data width as parameters
`define ADDR_WIDTH 16   // 16-bit address width
`define DATA_WIDTH 32   // 32-bit data width

// Optionally define other system-wide parameters
`define CLOCK_FREQ 100   // Clock frequency in MHz
`define RESET_ACTIVE_LOW 1   // 1 for active-low reset
